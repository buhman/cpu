`define BASE_SRC_RS1 1'b0
`define BASE_SRC_PC  1'b1

`define COND_NEVER 2'd0
`define COND_ALWAYS 2'd1
`define COND_EQ_ZERO 2'd2
`define COND_NEQ_ZERO 2'd3
