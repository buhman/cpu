`define ENCDEC_ZERO 2'b00
`define ENCDEC_BYTE 2'b01
`define ENCDEC_HALF 2'b10
`define ENCDEC_WORD 2'b11
