`ifdef VERILATOR
`define IMEM_INIT_PATH "../../aoc2020/day12/part1.imem"
`define DMEM_INIT_PATH "../../aoc2020/day12/input.dmem"
`else
`define IMEM_INIT_PATH "test/mret.imem"
`define DMEM_INIT_PATH "test/mret.imem"
`endif
