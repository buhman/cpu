`define ALU_A_ZERO 2'd0
`define ALU_A_PC   2'd1
`define ALU_A_RS1  2'd2

`define ALU_B_IMM  1'd0
`define ALU_B_RS2  1'd1
