`define RD_SRC_ALU_Y      2'b00
`define RD_SRC_DMEM_RDATA 2'b01
`define RD_SRC_PC_4       2'b10
